--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:19:48 11/12/2018
-- Design Name:   
-- Module Name:   /home/msca8h/Projects/EEE3163-pcfg/counter_test.vhd
-- Project Name:  pcfg
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: counter
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

ENTITY counter_test IS
END counter_test;

ARCHITECTURE behavior OF counter_test IS 
  
  -- Component Declaration for the Unit Under Test (UUT)
  
  COMPONENT counter
    PORT(
      clk  : IN  std_logic;
      ce   : IN  std_logic;
      sclr : IN  std_logic;
      q    : OUT std_logic_vector(10 downto 0)
      );
  END COMPONENT;
  

  --Inputs
  signal clk  : std_logic := '0';
  signal ce   : std_logic := '0';
  signal sclr : std_logic := '0';

  --Outputs
  signal q : std_logic_vector (10 downto 0);

  -- Clock period definitions
  constant clk_period : time := 10 ns;
  
BEGIN
  
  -- Instantiate the Unit Under Test (UUT)
  uut: counter PORT MAP (
    clk  => clk,
    ce   => ce,
    sclr => sclr,
    q    => q
    );

  -- Clock process definitions
  clk_process :process
  begin
    clk <= '0';
    wait for clk_period/2;
    clk <= '1';
    wait for clk_period/2;
  end process;
  

  -- Stimulus process
  stim_proc: process
  begin		
    -- hold reset state for 100 ns.
    wait for 1 ns;	
    sclr <= '1';
    wait for 10 ns;	
    sclr <= '0';
    wait for clk_period * 2;	
    ce <= '1';
    wait for clk_period * 5;	
    ce <= '0';
    wait for clk_period * 5;	
    ce <= '1';
    wait for clk_period * 5;	
    ce <= '0';
    wait for clk_period * 5;	
    sclr <= '1';
    wait for clk_period;	
    sclr <= '0';
    wait for clk_period * 5;	
    ce <= '1';
    wait for clk_period * 5;	
    ce <= '0';

    -- insert stimulus here 

    wait;
  end process;

END;
